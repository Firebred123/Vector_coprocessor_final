// include/custom_opcodes.vh
`define OPCODE_CUSTOM0 7'b0001011
`define FUNCT7_VLD   7'b0000001
`define FUNCT7_VST   7'b0000010
`define FUNCT7_VMAC  7'b0000011
